//`define MDU_ENABLE 1