//`define MDU_ENABLE 1
//`define UNALIGNED_ENABLE 1
//`define CSR_ENABLE 1
//`define RV32E 1