`define UART_ENABLE 1
`define GPIO_ENABLE 1
`define LED_ENABLE  1